// by KK

`timescale 1 ns / 1 ps

module top (
    input  wire clk,
    input wire rst,
    input  wire rx,
    input  wire sendBtn,
    output logic tx,
    output logic [3:0] an,
    output logic [6:0] seg,
    output logic dp
);

endmodule
