/**
 * San Jose State University
 * EE178 Lab #4
 * Author: prof. Eric Crabilla
 *
 * Modified by:
 * 2023  AGH University of Science and Technology
 * MTM UEC2
 * Piotr Kaczmarczyk
 *
 * Description:
 * The project top module.
 */

`timescale 1 ns / 1 ps

module top_vga (
    input  logic clk,
    input  logic clk100MHz,
    input  logic rst,
    output logic vs,
    output logic hs,
    output logic [3:0] r,
    output logic [3:0] g,
    output logic [3:0] b,

    inout logic ps2_clk,
    inout logic ps2_data
);


/**
 * Local variables and signals
 */

// VGA signals from background timing, rect, and mouse
vga_if vga_tim(), vga_bg(), vga_rect(), vga_mouse();
/**
 * Signals assignments
 */

assign vs = vga_mouse.vsync;
assign hs = vga_mouse.hsync;
assign {r,g,b} = vga_mouse.rgb;

logic [11:0] xpos;
logic [11:0] ypos;
logic [11:0] xpos_nxt;
logic [11:0] ypos_nxt;

always_ff @(posedge clk) begin
    if(rst) begin
        xpos <= '0;
        ypos <= '0;
    end else begin
        xpos <= xpos_nxt;
        ypos <= ypos_nxt;
    end
end

/**
 * Submodules instances
 */

vga_timing u_vga_timing (
    .clk,
    .rst,
    .vga(vga_tim)
);

draw_bg u_draw_bg (
    .clk,
    .rst,

    .vga_in(vga_tim),
    .vga_out(vga_bg)
);

draw_rect u_draw_rect (
    .clk,
    .rst,

    .x(xpos),
    .y(ypos),

    .vga_in(vga_bg),
    .vga_out(vga_rect)
);

draw_mouse u_draw_mouse (
    .clk,
    .rst,

    .x(xpos),
    .y(ypos),
    
    .vga_in(vga_rect),
    .vga_out(vga_mouse)
);

MouseCtl u_MouseCtl (
    .clk(clk100MHz),
    .rst,
    .ps2_clk,
    .ps2_data,
    .xpos(xpos_nxt),
    .ypos(ypos_nxt),

    .zpos(),
    .value(),
    .left(),
    .middle(),
    .right(),
    .setx(),
    .sety(),
    .setmax_x(),
    .setmax_y(),
    .new_event()
);

endmodule
