// by KK

package commands_pkg;

localparam ADD  = 3'b000;
localparam SUB  = 3'b001;
localparam AND  = 3'b010;
localparam OR   = 3'b011;
localparam NOP  = 3'b111;
localparam LDA  = 3'b100;
localparam LDB  = 3'b101;

localparam B1   = 3'b010;
localparam BR   = 3'b010;
localparam BN0  = 3'b101;

endpackage