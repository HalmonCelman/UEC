/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Piotr Kaczmarczyk
 *
 * Description:
 * Package with vga related constants.
 */

package rect_pkg;

localparam RECT_WIDTH=48;
localparam RECT_HEIGHT=64;

endpackage
